-- megafunction wizard: %ALTPLL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altpll 

-- ============================================================
-- File Name: uda1380pll.vhd
-- Megafunction Name(s):
-- 			altpll
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Full Version
-- ************************************************************

--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.

library ieee;
use ieee.std_logic_1164.all;

library altera_mf;
use altera_mf.all;

entity uda1380pll is
    port(
        inclk0 : in  std_logic := '0';
        c0     : out std_logic;
        locked : out std_logic);
end uda1380pll;

architecture SYN of uda1380pll is

    signal sub_wire0    : std_logic_vector(4 downto 0);
    signal sub_wire1    : std_logic;
    signal sub_wire2    : std_logic;
    signal sub_wire3    : std_logic;
    signal sub_wire4    : std_logic_vector(1 downto 0);
    signal sub_wire5_bv : BIT_VECTOR(0 downto 0);
    signal sub_wire5    : std_logic_vector(0 downto 0);

    component altpll
        generic(
            bandwidth_type          : string;
            clk0_divide_by          : NATURAL;
            clk0_duty_cycle         : NATURAL;
            clk0_multiply_by        : NATURAL;
            clk0_phase_shift        : string;
            compensate_clock        : string;
            inclk0_input_frequency  : NATURAL;
            intended_device_family  : string;
            lpm_hint                : string;
            lpm_type                : string;
            operation_mode          : string;
            pll_type                : string;
            port_activeclock        : string;
            port_areset             : string;
            port_clkbad0            : string;
            port_clkbad1            : string;
            port_clkloss            : string;
            port_clkswitch          : string;
            port_configupdate       : string;
            port_fbin               : string;
            port_inclk0             : string;
            port_inclk1             : string;
            port_locked             : string;
            port_pfdena             : string;
            port_phasecounterselect : string;
            port_phasedone          : string;
            port_phasestep          : string;
            port_phaseupdown        : string;
            port_pllena             : string;
            port_scanaclr           : string;
            port_scanclk            : string;
            port_scanclkena         : string;
            port_scandata           : string;
            port_scandataout        : string;
            port_scandone           : string;
            port_scanread           : string;
            port_scanwrite          : string;
            port_clk0               : string;
            port_clk1               : string;
            port_clk2               : string;
            port_clk3               : string;
            port_clk4               : string;
            port_clk5               : string;
            port_clkena0            : string;
            port_clkena1            : string;
            port_clkena2            : string;
            port_clkena3            : string;
            port_clkena4            : string;
            port_clkena5            : string;
            port_extclk0            : string;
            port_extclk1            : string;
            port_extclk2            : string;
            port_extclk3            : string;
            self_reset_on_loss_lock : string;
            width_clock             : NATURAL);
        port(
            clk    : out std_logic_vector(4 downto 0);
            inclk  : in  std_logic_vector(1 downto 0);
            locked : out std_logic);
    end component;

begin
    sub_wire5_bv(0 downto 0) <= "0";
    sub_wire5                <= To_stdlogicvector(sub_wire5_bv);
    sub_wire1                <= sub_wire0(0);
    c0                       <= sub_wire1;
    locked                   <= sub_wire2;
    sub_wire3                <= inclk0;
    sub_wire4                <= sub_wire5(0 downto 0) & sub_wire3;

    altpll_component : altpll
        generic map(
            bandwidth_type          => "AUTO",
            clk0_divide_by          => 3125,
            clk0_duty_cycle         => 50,
            clk0_multiply_by        => 768,
            clk0_phase_shift        => "0",
            compensate_clock        => "CLK0",
            inclk0_input_frequency  => 20000,
            intended_device_family  => "Cyclone IV E",
            lpm_hint                => "CBX_MODULE_PREFIX=uda1380pll",
            lpm_type                => "altpll",
            operation_mode          => "NORMAL",
            pll_type                => "AUTO",
            port_activeclock        => "PORT_UNUSED",
            port_areset             => "PORT_UNUSED",
            port_clkbad0            => "PORT_UNUSED",
            port_clkbad1            => "PORT_UNUSED",
            port_clkloss            => "PORT_UNUSED",
            port_clkswitch          => "PORT_UNUSED",
            port_configupdate       => "PORT_UNUSED",
            port_fbin               => "PORT_UNUSED",
            port_inclk0             => "PORT_USED",
            port_inclk1             => "PORT_UNUSED",
            port_locked             => "PORT_USED",
            port_pfdena             => "PORT_UNUSED",
            port_phasecounterselect => "PORT_UNUSED",
            port_phasedone          => "PORT_UNUSED",
            port_phasestep          => "PORT_UNUSED",
            port_phaseupdown        => "PORT_UNUSED",
            port_pllena             => "PORT_UNUSED",
            port_scanaclr           => "PORT_UNUSED",
            port_scanclk            => "PORT_UNUSED",
            port_scanclkena         => "PORT_UNUSED",
            port_scandata           => "PORT_UNUSED",
            port_scandataout        => "PORT_UNUSED",
            port_scandone           => "PORT_UNUSED",
            port_scanread           => "PORT_UNUSED",
            port_scanwrite          => "PORT_UNUSED",
            port_clk0               => "PORT_USED",
            port_clk1               => "PORT_UNUSED",
            port_clk2               => "PORT_UNUSED",
            port_clk3               => "PORT_UNUSED",
            port_clk4               => "PORT_UNUSED",
            port_clk5               => "PORT_UNUSED",
            port_clkena0            => "PORT_UNUSED",
            port_clkena1            => "PORT_UNUSED",
            port_clkena2            => "PORT_UNUSED",
            port_clkena3            => "PORT_UNUSED",
            port_clkena4            => "PORT_UNUSED",
            port_clkena5            => "PORT_UNUSED",
            port_extclk0            => "PORT_UNUSED",
            port_extclk1            => "PORT_UNUSED",
            port_extclk2            => "PORT_UNUSED",
            port_extclk3            => "PORT_UNUSED",
            self_reset_on_loss_lock => "OFF",
            width_clock             => 5)
        port map(
            inclk  => sub_wire4,
            clk    => sub_wire0,
            locked => sub_wire2);

end SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ACTIVECLK_CHECK string "0"
-- Retrieval info: PRIVATE: BANDWIDTH string "1.000"
-- Retrieval info: PRIVATE: BANDWIDTH_FEATURE_ENABLED string "1"
-- Retrieval info: PRIVATE: BANDWIDTH_FREQ_UNIT string "MHz"
-- Retrieval info: PRIVATE: BANDWIDTH_PRESET string "Low"
-- Retrieval info: PRIVATE: BANDWIDTH_USE_AUTO string "1"
-- Retrieval info: PRIVATE: BANDWIDTH_USE_PRESET string "0"
-- Retrieval info: PRIVATE: CLKBAD_SWITCHOVER_CHECK string "0"
-- Retrieval info: PRIVATE: CLKLOSS_CHECK string "0"
-- Retrieval info: PRIVATE: CLKSWITCH_CHECK string "0"
-- Retrieval info: PRIVATE: CNX_NO_COMPENSATE_RADIO string "0"
-- Retrieval info: PRIVATE: CREATE_CLKBAD_CHECK string "0"
-- Retrieval info: PRIVATE: CREATE_INCLK1_CHECK string "0"
-- Retrieval info: PRIVATE: CUR_DEDICATED_CLK string "c0"
-- Retrieval info: PRIVATE: CUR_FBIN_CLK string "c0"
-- Retrieval info: PRIVATE: DEVICE_SPEED_GRADE string "8"
-- Retrieval info: PRIVATE: DIV_FACTOR0 NUMERIC "297"
-- Retrieval info: PRIVATE: DUTY_CYCLE0 string "50.00000000"
-- Retrieval info: PRIVATE: EFF_OUTPUT_FREQ_VALUE0 string "12.288000"
-- Retrieval info: PRIVATE: EXPLICIT_SWITCHOVER_COUNTER string "0"
-- Retrieval info: PRIVATE: EXT_FEEDBACK_RADIO string "0"
-- Retrieval info: PRIVATE: GLOCKED_COUNTER_EDIT_CHANGED string "1"
-- Retrieval info: PRIVATE: GLOCKED_FEATURE_ENABLED string "0"
-- Retrieval info: PRIVATE: GLOCKED_MODE_CHECK string "0"
-- Retrieval info: PRIVATE: GLOCK_COUNTER_EDIT NUMERIC "1048575"
-- Retrieval info: PRIVATE: HAS_MANUAL_SWITCHOVER string "1"
-- Retrieval info: PRIVATE: INCLK0_FREQ_EDIT string "50.000"
-- Retrieval info: PRIVATE: INCLK0_FREQ_UNIT_COMBO string "MHz"
-- Retrieval info: PRIVATE: INCLK1_FREQ_EDIT string "100.000"
-- Retrieval info: PRIVATE: INCLK1_FREQ_EDIT_CHANGED string "1"
-- Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_CHANGED string "1"
-- Retrieval info: PRIVATE: INCLK1_FREQ_UNIT_COMBO string "MHz"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY string "Cyclone IV E"
-- Retrieval info: PRIVATE: INT_FEEDBACK__MODE_RADIO string "1"
-- Retrieval info: PRIVATE: LOCKED_OUTPUT_CHECK string "1"
-- Retrieval info: PRIVATE: LONG_SCAN_RADIO string "1"
-- Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE string "Not Available"
-- Retrieval info: PRIVATE: LVDS_MODE_DATA_RATE_DIRTY NUMERIC "0"
-- Retrieval info: PRIVATE: LVDS_PHASE_SHIFT_UNIT0 string "deg"
-- Retrieval info: PRIVATE: MIG_DEVICE_SPEED_GRADE string "Any"
-- Retrieval info: PRIVATE: MIRROR_CLK0 string "0"
-- Retrieval info: PRIVATE: MULT_FACTOR0 NUMERIC "73"
-- Retrieval info: PRIVATE: NORMAL_MODE_RADIO string "1"
-- Retrieval info: PRIVATE: OUTPUT_FREQ0 string "12.28800000"
-- Retrieval info: PRIVATE: OUTPUT_FREQ_MODE0 string "1"
-- Retrieval info: PRIVATE: OUTPUT_FREQ_UNIT0 string "MHz"
-- Retrieval info: PRIVATE: PHASE_RECONFIG_FEATURE_ENABLED string "1"
-- Retrieval info: PRIVATE: PHASE_RECONFIG_INPUTS_CHECK string "0"
-- Retrieval info: PRIVATE: PHASE_SHIFT0 string "0.00000000"
-- Retrieval info: PRIVATE: PHASE_SHIFT_STEP_ENABLED_CHECK string "0"
-- Retrieval info: PRIVATE: PHASE_SHIFT_UNIT0 string "deg"
-- Retrieval info: PRIVATE: PLL_ADVANCED_PARAM_CHECK string "0"
-- Retrieval info: PRIVATE: PLL_ARESET_CHECK string "0"
-- Retrieval info: PRIVATE: PLL_AUTOPLL_CHECK NUMERIC "1"
-- Retrieval info: PRIVATE: PLL_ENHPLL_CHECK NUMERIC "0"
-- Retrieval info: PRIVATE: PLL_FASTPLL_CHECK NUMERIC "0"
-- Retrieval info: PRIVATE: PLL_FBMIMIC_CHECK string "0"
-- Retrieval info: PRIVATE: PLL_LVDS_PLL_CHECK NUMERIC "0"
-- Retrieval info: PRIVATE: PLL_PFDENA_CHECK string "0"
-- Retrieval info: PRIVATE: PLL_TARGET_HARCOPY_CHECK NUMERIC "0"
-- Retrieval info: PRIVATE: PRIMARY_CLK_COMBO string "inclk0"
-- Retrieval info: PRIVATE: RECONFIG_FILE string "uda1380pll.mif"
-- Retrieval info: PRIVATE: SACN_INPUTS_CHECK string "0"
-- Retrieval info: PRIVATE: SCAN_FEATURE_ENABLED string "1"
-- Retrieval info: PRIVATE: SELF_RESET_LOCK_LOSS string "0"
-- Retrieval info: PRIVATE: SHORT_SCAN_RADIO string "0"
-- Retrieval info: PRIVATE: SPREAD_FEATURE_ENABLED string "0"
-- Retrieval info: PRIVATE: SPREAD_FREQ string "50.000"
-- Retrieval info: PRIVATE: SPREAD_FREQ_UNIT string "KHz"
-- Retrieval info: PRIVATE: SPREAD_PERCENT string "0.500"
-- Retrieval info: PRIVATE: SPREAD_USE string "0"
-- Retrieval info: PRIVATE: SRC_SYNCH_COMP_RADIO string "0"
-- Retrieval info: PRIVATE: STICKY_CLK0 string "1"
-- Retrieval info: PRIVATE: SWITCHOVER_COUNT_EDIT NUMERIC "1"
-- Retrieval info: PRIVATE: SWITCHOVER_FEATURE_ENABLED string "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX string "0"
-- Retrieval info: PRIVATE: USE_CLK0 string "1"
-- Retrieval info: PRIVATE: USE_CLKENA0 string "0"
-- Retrieval info: PRIVATE: USE_MIL_SPEED_GRADE NUMERIC "0"
-- Retrieval info: PRIVATE: ZERO_DELAY_RADIO string "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: BANDWIDTH_TYPE string "AUTO"
-- Retrieval info: CONSTANT: CLK0_DIVIDE_BY NUMERIC "3125"
-- Retrieval info: CONSTANT: CLK0_DUTY_CYCLE NUMERIC "50"
-- Retrieval info: CONSTANT: CLK0_MULTIPLY_BY NUMERIC "768"
-- Retrieval info: CONSTANT: CLK0_PHASE_SHIFT string "0"
-- Retrieval info: CONSTANT: COMPENSATE_CLOCK string "CLK0"
-- Retrieval info: CONSTANT: INCLK0_INPUT_FREQUENCY NUMERIC "20000"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY string "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_TYPE string "altpll"
-- Retrieval info: CONSTANT: OPERATION_MODE string "NORMAL"
-- Retrieval info: CONSTANT: PLL_TYPE string "AUTO"
-- Retrieval info: CONSTANT: PORT_ACTIVECLOCK string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ARESET string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_CLKBAD0 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_CLKBAD1 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_CLKLOSS string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_CLKSWITCH string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_CONFIGUPDATE string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FBIN string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_INCLK0 string "PORT_USED"
-- Retrieval info: CONSTANT: PORT_INCLK1 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_LOCKED string "PORT_USED"
-- Retrieval info: CONSTANT: PORT_PFDENA string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_PHASECOUNTERSELECT string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_PHASEDONE string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_PHASESTEP string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_PHASEUPDOWN string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_PLLENA string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANACLR string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANCLK string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANCLKENA string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANDATA string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANDATAOUT string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANDONE string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANREAD string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SCANWRITE string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clk0 string "PORT_USED"
-- Retrieval info: CONSTANT: PORT_clk1 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clk2 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clk3 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clk4 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clk5 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clkena0 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clkena1 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clkena2 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clkena3 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clkena4 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_clkena5 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_extclk0 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_extclk1 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_extclk2 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_extclk3 string "PORT_UNUSED"
-- Retrieval info: CONSTANT: SELF_RESET_ON_LOSS_LOCK string "OFF"
-- Retrieval info: CONSTANT: WIDTH_CLOCK NUMERIC "5"
-- Retrieval info: USED_PORT: @clk 0 0 5 0 OUTPUT_CLK_EXT VCC "@clk[4..0]"
-- Retrieval info: USED_PORT: @inclk 0 0 2 0 INPUT_CLK_EXT VCC "@inclk[1..0]"
-- Retrieval info: USED_PORT: c0 0 0 0 0 OUTPUT_CLK_EXT VCC "c0"
-- Retrieval info: USED_PORT: inclk0 0 0 0 0 INPUT_CLK_EXT GND "inclk0"
-- Retrieval info: USED_PORT: locked 0 0 0 0 OUTPUT GND "locked"
-- Retrieval info: CONNECT: @inclk 0 0 1 1 GND 0 0 0 0
-- Retrieval info: CONNECT: @inclk 0 0 1 0 inclk0 0 0 0 0
-- Retrieval info: CONNECT: c0 0 0 0 0 @clk 0 0 1 0
-- Retrieval info: CONNECT: locked 0 0 0 0 @locked 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL uda1380pll.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL uda1380pll.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL uda1380pll.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL uda1380pll.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL uda1380pll.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL uda1380pll_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: CBX_MODULE_PREFIX: ON
